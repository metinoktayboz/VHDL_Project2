----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:43:00 11/10/2019 
-- Design Name: 
-- Module Name:    NotA - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity NotA is
Port(
 a1 : in STD_LOGIC_VECTOR(3 downto 0);
out1: out STD_LOGIC_VECTOR(3 downto 0)
);end NotA;

architecture Behavioral of NotA is

begin
out1 <= (not a1);


end Behavioral;


